package fifopkg;

  `include "rstgen.sv"
  `include "write_readtest.sv"
  `include "underflow_test.sv"
  `include "overflow_test.sv"
  `include "empty_test.sv"
  `include "full_test.sv"
  `include "result.sv"
  `include "reset_test.sv"
  `include "runtest.sv"
  
endpackage

